
entity multiplexer is
	port(a,b,c,d, sel1, sel2: in bit;
	    y: out bit);
end entity;

architecture behavior of multiplexer is
begin
	
end architecture;
